<svg width="34" height="31" viewBox="0 0 34 31" fill="none" xmlns="http://www.w3.org/2000/svg">
<g opacity="0.5">
<path d="M20 15.5393L14.75 19.3101V11.7684L20 15.5393Z" fill="black" stroke="black" stroke-width="2.74646" stroke-linecap="round" stroke-linejoin="round"/>
<path d="M2 16.8732V14.2052C2 8.74619 2 6.01674 3.35823 4.26053C4.71648 2.50431 6.85484 2.42829 11.1315 2.27625C13.1581 2.20421 15.2282 2.15259 17 2.15259C18.7718 2.15259 20.842 2.20421 22.8685 2.27625C27.1451 2.42829 29.2835 2.50431 30.6417 4.26053C32 6.01674 32 8.74619 32 14.2052V16.8732C32 22.3321 32 25.0616 30.6417 26.8177C29.2835 28.574 27.1453 28.6499 22.8686 28.8021C20.842 28.8741 18.7718 28.9258 17 28.9258C15.2282 28.9258 13.158 28.8741 11.1314 28.8021C6.85476 28.6499 4.71645 28.574 3.35822 26.8177C2 25.0616 2 22.3321 2 16.8732Z" stroke="black" stroke-width="2.74646"/>
</g>
</svg>
